** Profile: "SCHEMATIC1-Workshop"  [ C:\USERS\AMMAR ISSA\DESKTOP\Workshop\workshop-SCHEMATIC1-Workshop.sim ] 

** Creating circuit file "workshop-SCHEMATIC1-Workshop.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5ms 0 0.1ms SKIPBP 
.OPTIONS DIGINITSTATE= 1
.OPTIONS DIGIOLVL= 2
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\workshop-SCHEMATIC1.net" 


.END
